library ieee;
use ieee.std_logic_1164.all;

entity ss7 is
port
	(
	bcd : in std_logic_vector(3 downto 0); --Recibe un numero entero como entrada.
	HEX : out std_logic_vector(6 downto 0) --Tiene un arreglo de 7 bits como salida.
	);
end entity;

architecture a of ss7 is
begin
	with bcd select
	HEX <= 
		"1000000" when "0000",
		"1111001" when "0001",
		"0100100" when "0010",
		"0110000" when "0011",
		"0011001" when "0100",
		"0010010" when "0101",
		"0000010" when "0110",
		"1111000" when "0111",
		"0000000" when "1000",
		"0011000" when "1001",
	   "0000000" when others;	--Solo se tomarán en cuenta enteros de 0 a 9.
end architecture;
